counter_30_inst : counter_30 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
