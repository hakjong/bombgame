counter_16_inst : counter_16 PORT MAP (
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
