counter_48mhz_inst : counter_48mhz PORT MAP (
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
